module

endmodule